module MyOperators( // @[:@3.2]
  input        clock, // @[:@4.4]
  input        reset, // @[:@5.4]
  input  [3:0] io_in, // @[:@6.4]
  output [3:0] io_out_add, // @[:@6.4]
  output [3:0] io_out_sub, // @[:@6.4]
  output [3:0] io_out_mul // @[:@6.4]
);
  wire [3:0] _T_15; // @[ChiselBootcamp22.scala 22:23:@8.4]
  wire [2:0] _T_16; // @[ChiselBootcamp22.scala 22:23:@9.4]
  wire [2:0] _T_19; // @[ChiselBootcamp22.scala 23:23:@11.4]
  wire [2:0] _T_20; // @[ChiselBootcamp22.scala 23:23:@12.4]
  wire [1:0] _T_21; // @[ChiselBootcamp22.scala 23:23:@13.4]
  wire [4:0] _T_24; // @[ChiselBootcamp22.scala 24:23:@15.4]
  assign _T_15 = 3'h1 + 3'h4; // @[ChiselBootcamp22.scala 22:23:@8.4]
  assign _T_16 = _T_15[2:0]; // @[ChiselBootcamp22.scala 22:23:@9.4]
  assign _T_19 = 2'h2 - 2'h1; // @[ChiselBootcamp22.scala 23:23:@11.4]
  assign _T_20 = $unsigned(_T_19); // @[ChiselBootcamp22.scala 23:23:@12.4]
  assign _T_21 = _T_20[1:0]; // @[ChiselBootcamp22.scala 23:23:@13.4]
  assign _T_24 = 3'h4 * 3'h2; // @[ChiselBootcamp22.scala 24:23:@15.4]
  assign io_out_add = {{1'd0}, _T_16}; // @[ChiselBootcamp22.scala 22:16:@10.4]
  assign io_out_sub = {{2'd0}, _T_21}; // @[ChiselBootcamp22.scala 23:16:@14.4]
  assign io_out_mul = _T_24[3:0]; // @[ChiselBootcamp22.scala 24:16:@16.4]
endmodule
